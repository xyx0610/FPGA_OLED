module change_xy(
	input clk,
	input rst_n,
	input add_dec_x,
	input add_dec_y,
	output reg [6:0] x,
	output reg [5:0] y
);



endmodule